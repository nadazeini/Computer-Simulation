// Name: logic.v
// Module: 
// Input: 
// Output: 
//
// Notes: Common definitions
// 
//
// Revision History:
//
// Version	Date		Who		email			note
//------------------------------------------------------------------------------------------
//  1.0     Sep 02, 2014	Kaushik Patra	kpatra@sjsu.edu		Initial creation
//------------------------------------------------------------------------------------------
//
// 64-bit two's complement
module TWOSCOMP64(Y,A);
//output list
output [63:0] Y;
//input list
input [63:0] A;
wire [63:0] not_out;

wire null2;
genvar i;
generate
for(i=0;i<64;i=i+1)
begin : loop_2s_64
not not_inst(not_out[i],A[i]);
end
endgenerate
RC_ADD_SUB_64 adder(Y, null2 ,not_out, 64'b1, 1'b0);

endmodule

// 32-bit two's complement
module TWOSCOMP32(Y,A);
//output list
output [31:0] Y;
//input list
input [31:0] A;
wire [31:0] not_out;
//add wires
wire null1;
genvar j;
generate
for(j=0;j<32;j=j+1)
begin : loop_2s_32
not not_inst(not_out[j],A[j]);
end
endgenerate
RC_ADD_SUB_32 adder(Y, null1 ,not_out, 32'b1, 1'b0);
endmodule

//special registers
module REG32_PP(Q, D,LOAD, CLK, RESET);
	input CLK,LOAD,RESET;
	input [31:0] D;
	output [31:0] Q;
	wire [31:0] Qbar;
	//wire notR;
	parameter PATTERN = 32'h00000000;
	genvar i;
	generate
		for (i=0; i<32; i=i+1) begin : bitreg_gen_loop
			//not n(notR, RESET);
if(PATTERN[i]==0)
			REG1 r(.Q(Q[i]), .Qbar(Qbar), .nR(RESET), .D(D[i]), .L(LOAD), .C(CLK), .nP(1'b1));
else REG1 r(.Q(Q[i]), .Qbar(Qbar), .nR(1'b1), .D(D[i]), .L(LOAD), .C(CLK), .nP(RESET));
		end
	endgenerate

endmodule


// 32-bit registere +ve edge, Reset on RESET=0
module REG32(Q, D,LOAD, CLK, RESET);
	input CLK,LOAD,RESET;
	input [31:0] D;
	output [31:0] Q;
	wire Qbar;
	wire notR;
	
	genvar i;
	generate
		for (i=0; i<32; i=i+1) begin : bitreg_gen_loop
			//not n(notR, RESET);
			REG1 r(.Q(Q[i]), .Qbar(Qbar), .nR(1'b1), .D(D[i]), .L(LOAD), .C(CLK), .nP(RESET));
		end
	endgenerate

endmodule
// 1 bit register +ve edge, 
// Preset on nP=0, nR=1, reset on nP=1, nR=0;
// Undefined nP=0, nR=0
// normal operation nP=1, nR=1
module REG1(Q, Qbar, D, L, C, nP, nR);
	input nR, D, L, C, nP;
	output Q, Qbar;
	wire muxOut;
	wire flopOut;	
	 MUX1_2x1 m(muxOut, ff_out, D, L);

	D_FF b(.Q(ff_out), .Qbar(Qbar), .nR(nR), .D(muxOut), .C(C), .nP(nP));
	buf(Q, ff_out);
endmodule
// 1 bit flipflop +ve edge, 
// Preset on nP=0, nR=1, reset on nP=1, nR=0;
// Undefined nP=0, nR=0
// normal operation nP=1, nR=1
module D_FF(Q, Qbar, D, C,nP, nR);
	input nR, D, C, nP;
	output Q, Qbar;
	wire notD, notC, dout1, dout2;
D_LATCH dl(.Q(dout1), .Qbar(dout2), .D(D), .C(C), .nP(nP), .nR(nR));
SR_LATCH srl(.Q(Q),.Qbar(Qbar),.S(dout1),.R(dout2),.C(C),.nP(nP),.nR(nR));
endmodule

// 1 bit D latch
// Preset on nP=0, nR=1, reset on nP=1, nR=0;
// Undefined nP=0, nR=0
// normal operation nP=1, nR=1
module D_LATCH(Q, Qbar, D, C, nP, nR);
input D, C;
input nP, nR;
output Q,Qbar;
wire Dbar;


wire Y,Ybar;
wire [9:0] out;
wire dOut1,dOut2;
	not invD(notD, D);
not invC(notC, C);
	nand nand1(out[2], D, notC);
	nand nand2(out[3], notD, notC);
	nand nand3(dOut1, nR, out[2], dOut2);
	nand nand4(dOut2, dOut1, out[3], nP);
buf b1(Q, dOut1);
buf b2(Qbar, dOut2);
endmodule
// 1 bit SR latch
// Preset on nP=0, nR=1, reset on nP=1, nR=0;
// Undefined nP=0, nR=0
// normal operation nP=1, nR=1
module SR_LATCH(Q,Qbar,S,R,C,nP,nR);
input S,R,C;
input nP, nR;
output Q,Qbar;
wire out[9:0];
	not invC(notC, C);
	nand nand1(out[6], S, C);
	nand nand2(out[7], C, R);
	nand nand3(out[8], nR, out[6], out[9]);
	nand nand4(out[9], out[8], out[7], nP);
	buf bufQ(Q, out[8]);
	buf bufQbar(Qbar, out[9]);
endmodule


// 5x32 Line decoder
module DECODER_5x32(D,I);
// output
output [31:0] D;
// input
input [4:0] I;

wire [16:0]d; //half of 32 //delete this
 DECODER_4x16 d4x16(d[15:0],I[3:0]);
not not_inst(d[16],I[4]);
genvar i;
generate
for(i=0;i<16;i=i+1)
begin :d_loop
and and1(D[i],d[i],d[16]);
and and2(D[i+16],I[4],d[i]);
end
endgenerate
endmodule

// 4x16 Line decoder
module DECODER_4x16(D,I);
// output
output [15:0] D;
// input
input [3:0] I;
wire [8:0]d;
 DECODER_3x8 d3x8(d[7:0],I[2:0]);
not not_inst(d[8],I[3]);
genvar i;
generate
for(i=0;i<8;i=i+1)
begin :d_loop
and and1(D[i],d[i],d[8]);
and and2(D[i+8],I[3],d[i]);
end
endgenerate


endmodule

// 3x8 Line decoder
module DECODER_3x8(D,I);
// output
output [7:0] D;
// input
input [2:0] I;
wire [4:0]d;
DECODER_2x4 d2x4(d[3:0],I[1:0]); //leave one out for third input
not inst(d[4],I[2]);
//use generate cause faster
genvar i;
generate
for(i=0;i<4;i=i+1) 
begin : decoder_loop
and and1(D[i],d[4],d[i]);
and and2(D[i+4],I[2],d[i]);
end
endgenerate
endmodule

// 2x4 Line decoder
module DECODER_2x4(D,I);
// output
output [3:0] D;
// input
input [1:0] I;

wire W[1:0];

not not1(W[0],I[0]);//first inverter
not not2(W[1],I[1]);//second inverter
and and1(D[0],W[0],W[1]);
and and2(D[1],W[1],I[0]);
and and3(D[2],W[0],I[1]);
and and4(D[3],I[0],I[1]);


endmodule




//implement 3 input NAND
module NAND_3 (out,A,B,C);


input A,B,C;
output out;
wire out_wire[1:0];
and and_inst(out_wire[0],A,B);
and and1 (out_wire[1],out_wire[0],C);
not not_inst(out,out_wire[1]);
endmodule












                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  
`timescale 1ns/1ps
module mux_tb;
/*reg S,I0, I1;
wire Y;
//testing 1 bit mux 2 by 1
MUX1_2x1 mux1_2x1(.Y(Y),.I0(I0),.I1(I1),.S(S));
initial 
begin
#5 $write("\n Testing 1 bit mux 2x1 \n");
#5 S=0; I0=0; I1=0;
#5 $write("\n control is:%d I0=%d I1=%d result is:%d\n",S,I0,I1,Y);
#5 S=0; I0=1; I1=0;
#5 $write("\n control is:%d I0=%d I1=%d result is:%d\n",S,I0,I1,Y);
#5 S=0; I0=0; I1=1;
#5 $write("\n control is:%d I0=%d I1=%d result is:%d\n",S,I0,I1,Y);
#5 S=0; I0=1; I1=1;
#5 $write("\n control is:%d I0=%d I1=%d result is:%d\n",S,I0,I1,Y);
#5 S=1; I0=0; I1=0;
#5 $write("\n control is:%d I0=%d I1=%d result is:%d\n",S,I0,I1,Y);
#5 S=1; I0=1; I1=0;
#5 $write("\n control is:%d I0=%d I1=%d result is:%d\n",S,I0,I1,Y);
#5 S=1; I0=0; I1=1;
#5 $write("\n control is:%d I0=%d I1=%d result is:%d\n",S,I0,I1,Y);
#5 S=1; I0=1; I1=1;
#5 $write("\n control is:%d I0=%d I1=%d result is:%d\n",S,I0,I1,Y);
end */


//TEST FOR 2x1 MUX
/*reg [31:0] I0, I1;
reg S;
wire [31:0] Y;
MUX32_2x1 mux32_2x1(.Y(Y),.I0(I0),.I1(I1),.S(S));
initial 
begin
#5 $write("\n Testing 32 bit mux 2x1 \n");
#5 S=0; I0=0; I1=0;
#5 $write("\n control is:%d I0=%d I1=%d result is:%d\n",S,I0,I1,Y);
#5 S=0; I0=1; I1=0;
#5 $write("\n control is:%d I0=%d I1=%d result is:%d\n",S,I0,I1,Y);
#5 S=0; I0=0; I1=1;
#5 $write("\n control is:%d I0=%d I1=%d result is:%d\n",S,I0,I1,Y);
#5 S=0; I0=1; I1=1;
#5 $write("\n control is:%d I0=%d I1=%d result is:%d\n",S,I0,I1,Y);
#5 S=1; I0=0; I1=0;
#5 $write("\n control is:%d I0=%d I1=%d result is:%d\n",S,I0,I1,Y);
#5 S=1; I0=1; I1=0;
#5 $write("\n control is:%d I0=%d I1=%d result is:%d\n",S,I0,I1,Y);
#5 S=1; I0=0; I1=1;
#5 $write("\n control is:%d I0=%d I1=%d result is:%d\n",S,I0,I1,Y);
#5 S=1; I0=1; I1=1;
#5 $write("\n control is:%d I0=%d I1=%d result is:%d\n",S,I0,I1,Y);
end
endmodule */

//TEST FOR 4x1 MUX
/*reg [31:0] I0, I1,I2,I3;
reg [1:0] S;
wire [31:0] Y,mux1out,mux2out;
MUX32_4x1 mux32_4x1(.Y(Y), .I0(I0), .I1(I1), .I2(I2), .I3(I3), .S(S));
initial 
begin
#5 $write("\n Testing 32 bit mux 4x1 \n");
#5 S=2'b00; I0=0; I1=1; I2=2; I3=3;
#5 $write(" control is:%b I0=%d I1=%d I2=%d I3=%d result is:%d\n",S,I0,I1,I2,I3,Y);
#5 S=2'b01; I0=0; I1=1; I2=2; I3=3;
#5 $write(" control is:%b I0=%d I1=%d I2=%d I3=%d result is:%d\n",S,I0,I1,I2,I3,Y);
#5 S=2'b10; I0=0; I1=1; I2=2; I3=3;
#5 $write(" control is:%b I0=%d I1=%d I2=%d I3=%d result is:%d\n",S,I0,I1,I2,I3,Y);
#5 S=2'b11; I0=0; I1=1; I2=2; I3=3;
#5 $write(" control is:%b I0=%d I1=%d I2=%d I3=%d result is:%d\n",S,I0,I1,I2,I3,Y);


end
endmodule 
*/


//TEST FOR 32x1 MUX

reg [31:0]  I0, I1, I2, I3, I4, I5, I6, I7;
reg [31:0] I8, I9, I10, I11, I12, I13, I14, I15;
reg [31:0] I16, I17, I18, I19, I20, I21, I22, I23;
reg [31:0] I24, I25, I26, I27, I28, I29, I30, I31;
reg [4:0] S;
wire [31:0] Y, mux16x1_out1,mux16x1_out2;
MUX32_32x1 mux32x1(.Y(Y),.I0(I0),.I1(I1),.I2(I2),.I3(I3),.I4(I4),.I5(I5),.I6(I6),.I7(I7),
.I8(I8),.I9(I9),.I10(I10),.I11(I11),.I12(I12),.I13(I13),.I14(I14),.I15(I15),.I16(I16),.I17(I17),.I18(I18),.I19(I19),.I20(I20),.I21(I21),
.I22(I22),.I23(I23),.I24(I24),.I25(I25),.I26(I26),.I27(I27),.I28(I28),.I29(I29),.I30(I30),
.I31(I31),.S(S));
initial
begin
#5 $write("\n Testing 32 bit mux 32x1 \n");
#5 S=5'b00000; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b I0=%d I1=%d I2=%d I3=%d I4=%d I5=%d I6=%d I7=%d
                     I8=%d, I9=%d I10=%d, I11=%d, I12=%d I13=%d I14=%d I15=%d
                     I16=%d I17=%d I18=%d I19=%d I20=%d I21=%d I22=%d I23=%d
                     I2=%d I25=%d I26=%d I27=%d I28=%d I29=%d I30=%d I31=%d result is:%d\n",S, I0, I1, I2, I3, I4, I5, I6, I7,
                     I8, I9, I10, I11, I12, I13, I14, I15,
                     I16, I17, I18, I19, I20, I21, I22, I23,
                     I24, I25, I26, I27, I28, I29, I30, I31,Y);
#5 S=5'b00001; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b00010; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b00011; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b00100; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b00101; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b00110; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b00111; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b01000; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b01001; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b01010; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b01011; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b01100; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b01101; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b01110; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b01111; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b10000; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b10001; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b10010; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b10011; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b10100; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b10101; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b10110; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b10111; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b11000; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b11001; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b11010; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b11011; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b11100; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b11101; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b11110; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
#5 S=5'b11111; I0=0; I1=1; I2=2;I3=3;I4=4;I5=5;I6=6;I7=7;I8=8;I9=9;I10=10;I11=11;
		I12=12;I13=13;I14=14;I15=15;I16=16;I17=17;I18=18;I19=19;I20=20;I21=21;
		I22=22;I23=23;I24=24;I25=25;I26=26;I27=27;I28=28;I29=29;I30=30;I31=31;
#5 $write("control is:%b result is:%d\n",S,Y);
end

endmodule 



